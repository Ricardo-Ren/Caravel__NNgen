magic
tech sky130A
magscale 1 2
timestamp 1654242109
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 290 1232 118864 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2410 119200 2466 120000
rect 3422 119200 3478 120000
rect 4434 119200 4490 120000
rect 5446 119200 5502 120000
rect 6458 119200 6514 120000
rect 7470 119200 7526 120000
rect 8482 119200 8538 120000
rect 9494 119200 9550 120000
rect 10506 119200 10562 120000
rect 11518 119200 11574 120000
rect 12530 119200 12586 120000
rect 13542 119200 13598 120000
rect 14554 119200 14610 120000
rect 15566 119200 15622 120000
rect 16578 119200 16634 120000
rect 17590 119200 17646 120000
rect 18602 119200 18658 120000
rect 19614 119200 19670 120000
rect 20626 119200 20682 120000
rect 21638 119200 21694 120000
rect 22650 119200 22706 120000
rect 23662 119200 23718 120000
rect 24582 119200 24638 120000
rect 25594 119200 25650 120000
rect 26606 119200 26662 120000
rect 27618 119200 27674 120000
rect 28630 119200 28686 120000
rect 29642 119200 29698 120000
rect 30654 119200 30710 120000
rect 31666 119200 31722 120000
rect 32678 119200 32734 120000
rect 33690 119200 33746 120000
rect 34702 119200 34758 120000
rect 35714 119200 35770 120000
rect 36726 119200 36782 120000
rect 37738 119200 37794 120000
rect 38750 119200 38806 120000
rect 39762 119200 39818 120000
rect 40774 119200 40830 120000
rect 41786 119200 41842 120000
rect 42798 119200 42854 120000
rect 43810 119200 43866 120000
rect 44822 119200 44878 120000
rect 45834 119200 45890 120000
rect 46846 119200 46902 120000
rect 47858 119200 47914 120000
rect 48778 119200 48834 120000
rect 49790 119200 49846 120000
rect 50802 119200 50858 120000
rect 51814 119200 51870 120000
rect 52826 119200 52882 120000
rect 53838 119200 53894 120000
rect 54850 119200 54906 120000
rect 55862 119200 55918 120000
rect 56874 119200 56930 120000
rect 57886 119200 57942 120000
rect 58898 119200 58954 120000
rect 59910 119200 59966 120000
rect 60922 119200 60978 120000
rect 61934 119200 61990 120000
rect 62946 119200 63002 120000
rect 63958 119200 64014 120000
rect 64970 119200 65026 120000
rect 65982 119200 66038 120000
rect 66994 119200 67050 120000
rect 68006 119200 68062 120000
rect 69018 119200 69074 120000
rect 70030 119200 70086 120000
rect 71042 119200 71098 120000
rect 72054 119200 72110 120000
rect 72974 119200 73030 120000
rect 73986 119200 74042 120000
rect 74998 119200 75054 120000
rect 76010 119200 76066 120000
rect 77022 119200 77078 120000
rect 78034 119200 78090 120000
rect 79046 119200 79102 120000
rect 80058 119200 80114 120000
rect 81070 119200 81126 120000
rect 82082 119200 82138 120000
rect 83094 119200 83150 120000
rect 84106 119200 84162 120000
rect 85118 119200 85174 120000
rect 86130 119200 86186 120000
rect 87142 119200 87198 120000
rect 88154 119200 88210 120000
rect 89166 119200 89222 120000
rect 90178 119200 90234 120000
rect 91190 119200 91246 120000
rect 92202 119200 92258 120000
rect 93214 119200 93270 120000
rect 94226 119200 94282 120000
rect 95238 119200 95294 120000
rect 96250 119200 96306 120000
rect 97170 119200 97226 120000
rect 98182 119200 98238 120000
rect 99194 119200 99250 120000
rect 100206 119200 100262 120000
rect 101218 119200 101274 120000
rect 102230 119200 102286 120000
rect 103242 119200 103298 120000
rect 104254 119200 104310 120000
rect 105266 119200 105322 120000
rect 106278 119200 106334 120000
rect 107290 119200 107346 120000
rect 108302 119200 108358 120000
rect 109314 119200 109370 120000
rect 110326 119200 110382 120000
rect 111338 119200 111394 120000
rect 112350 119200 112406 120000
rect 113362 119200 113418 120000
rect 114374 119200 114430 120000
rect 115386 119200 115442 120000
rect 116398 119200 116454 120000
rect 117410 119200 117466 120000
rect 118422 119200 118478 120000
rect 119434 119200 119490 120000
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60646 0 60702 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82266 0 82322 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87602 0 87658 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91466 0 91522 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103426 0 103482 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 105818 0 105874 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109498 0 109554 800
rect 109682 0 109738 800
rect 109958 0 110014 800
rect 110142 0 110198 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112074 0 112130 800
rect 112350 0 112406 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113822 0 113878 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115202 0 115258 800
rect 115478 0 115534 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116214 0 116270 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 116950 0 117006 800
rect 117134 0 117190 800
rect 117410 0 117466 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119802 0 119858 800
<< obsm2 >>
rect 110 119144 422 119354
rect 590 119144 1342 119354
rect 1510 119144 2354 119354
rect 2522 119144 3366 119354
rect 3534 119144 4378 119354
rect 4546 119144 5390 119354
rect 5558 119144 6402 119354
rect 6570 119144 7414 119354
rect 7582 119144 8426 119354
rect 8594 119144 9438 119354
rect 9606 119144 10450 119354
rect 10618 119144 11462 119354
rect 11630 119144 12474 119354
rect 12642 119144 13486 119354
rect 13654 119144 14498 119354
rect 14666 119144 15510 119354
rect 15678 119144 16522 119354
rect 16690 119144 17534 119354
rect 17702 119144 18546 119354
rect 18714 119144 19558 119354
rect 19726 119144 20570 119354
rect 20738 119144 21582 119354
rect 21750 119144 22594 119354
rect 22762 119144 23606 119354
rect 23774 119144 24526 119354
rect 24694 119144 25538 119354
rect 25706 119144 26550 119354
rect 26718 119144 27562 119354
rect 27730 119144 28574 119354
rect 28742 119144 29586 119354
rect 29754 119144 30598 119354
rect 30766 119144 31610 119354
rect 31778 119144 32622 119354
rect 32790 119144 33634 119354
rect 33802 119144 34646 119354
rect 34814 119144 35658 119354
rect 35826 119144 36670 119354
rect 36838 119144 37682 119354
rect 37850 119144 38694 119354
rect 38862 119144 39706 119354
rect 39874 119144 40718 119354
rect 40886 119144 41730 119354
rect 41898 119144 42742 119354
rect 42910 119144 43754 119354
rect 43922 119144 44766 119354
rect 44934 119144 45778 119354
rect 45946 119144 46790 119354
rect 46958 119144 47802 119354
rect 47970 119144 48722 119354
rect 48890 119144 49734 119354
rect 49902 119144 50746 119354
rect 50914 119144 51758 119354
rect 51926 119144 52770 119354
rect 52938 119144 53782 119354
rect 53950 119144 54794 119354
rect 54962 119144 55806 119354
rect 55974 119144 56818 119354
rect 56986 119144 57830 119354
rect 57998 119144 58842 119354
rect 59010 119144 59854 119354
rect 60022 119144 60866 119354
rect 61034 119144 61878 119354
rect 62046 119144 62890 119354
rect 63058 119144 63902 119354
rect 64070 119144 64914 119354
rect 65082 119144 65926 119354
rect 66094 119144 66938 119354
rect 67106 119144 67950 119354
rect 68118 119144 68962 119354
rect 69130 119144 69974 119354
rect 70142 119144 70986 119354
rect 71154 119144 71998 119354
rect 72166 119144 72918 119354
rect 73086 119144 73930 119354
rect 74098 119144 74942 119354
rect 75110 119144 75954 119354
rect 76122 119144 76966 119354
rect 77134 119144 77978 119354
rect 78146 119144 78990 119354
rect 79158 119144 80002 119354
rect 80170 119144 81014 119354
rect 81182 119144 82026 119354
rect 82194 119144 83038 119354
rect 83206 119144 84050 119354
rect 84218 119144 85062 119354
rect 85230 119144 86074 119354
rect 86242 119144 87086 119354
rect 87254 119144 88098 119354
rect 88266 119144 89110 119354
rect 89278 119144 90122 119354
rect 90290 119144 91134 119354
rect 91302 119144 92146 119354
rect 92314 119144 93158 119354
rect 93326 119144 94170 119354
rect 94338 119144 95182 119354
rect 95350 119144 96194 119354
rect 96362 119144 97114 119354
rect 97282 119144 98126 119354
rect 98294 119144 99138 119354
rect 99306 119144 100150 119354
rect 100318 119144 101162 119354
rect 101330 119144 102174 119354
rect 102342 119144 103186 119354
rect 103354 119144 104198 119354
rect 104366 119144 105210 119354
rect 105378 119144 106222 119354
rect 106390 119144 107234 119354
rect 107402 119144 108246 119354
rect 108414 119144 109258 119354
rect 109426 119144 110270 119354
rect 110438 119144 111282 119354
rect 111450 119144 112294 119354
rect 112462 119144 113306 119354
rect 113474 119144 114318 119354
rect 114486 119144 115330 119354
rect 115498 119144 116342 119354
rect 116510 119144 117354 119354
rect 117522 119144 118366 119354
rect 110 856 118478 119144
rect 222 800 238 856
rect 406 800 514 856
rect 682 800 698 856
rect 866 800 974 856
rect 1142 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1710 856
rect 1878 800 1894 856
rect 2062 800 2170 856
rect 2338 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2906 856
rect 3074 800 3090 856
rect 3258 800 3366 856
rect 3534 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4102 856
rect 4270 800 4378 856
rect 4546 800 4562 856
rect 4730 800 4838 856
rect 5006 800 5022 856
rect 5190 800 5298 856
rect 5466 800 5574 856
rect 5742 800 5758 856
rect 5926 800 6034 856
rect 6202 800 6218 856
rect 6386 800 6494 856
rect 6662 800 6770 856
rect 6938 800 6954 856
rect 7122 800 7230 856
rect 7398 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8426 856
rect 8594 800 8702 856
rect 8870 800 8886 856
rect 9054 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9622 856
rect 9790 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11094 856
rect 11262 800 11278 856
rect 11446 800 11554 856
rect 11722 800 11830 856
rect 11998 800 12014 856
rect 12182 800 12290 856
rect 12458 800 12474 856
rect 12642 800 12750 856
rect 12918 800 13026 856
rect 13194 800 13210 856
rect 13378 800 13486 856
rect 13654 800 13670 856
rect 13838 800 13946 856
rect 14114 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14682 856
rect 14850 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15418 856
rect 15586 800 15602 856
rect 15770 800 15878 856
rect 16046 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16614 856
rect 16782 800 16798 856
rect 16966 800 17074 856
rect 17242 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17810 856
rect 17978 800 17994 856
rect 18162 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18730 856
rect 18898 800 19006 856
rect 19174 800 19282 856
rect 19450 800 19466 856
rect 19634 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21398 856
rect 21566 800 21674 856
rect 21842 800 21858 856
rect 22026 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22870 856
rect 23038 800 23054 856
rect 23222 800 23330 856
rect 23498 800 23606 856
rect 23774 800 23790 856
rect 23958 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24526 856
rect 24694 800 24802 856
rect 24970 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26458 856
rect 26626 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27194 856
rect 27362 800 27378 856
rect 27546 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30782 856
rect 30950 800 31058 856
rect 31226 800 31242 856
rect 31410 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31978 856
rect 32146 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32714 856
rect 32882 800 32990 856
rect 33158 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35382 856
rect 35550 800 35566 856
rect 35734 800 35842 856
rect 36010 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36578 856
rect 36746 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37774 856
rect 37942 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38970 856
rect 39138 800 39154 856
rect 39322 800 39430 856
rect 39598 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40902 856
rect 41070 800 41086 856
rect 41254 800 41362 856
rect 41530 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42834 856
rect 43002 800 43018 856
rect 43186 800 43294 856
rect 43462 800 43478 856
rect 43646 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45686 856
rect 45854 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46882 856
rect 47050 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47618 856
rect 47786 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48538 856
rect 48706 800 48814 856
rect 48982 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49734 856
rect 49902 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50746 856
rect 50914 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51482 856
rect 51650 800 51666 856
rect 51834 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53138 856
rect 53306 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53874 856
rect 54042 800 54058 856
rect 54226 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55346 856
rect 55514 800 55530 856
rect 55698 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56266 856
rect 56434 800 56542 856
rect 56710 800 56726 856
rect 56894 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57462 856
rect 57630 800 57738 856
rect 57906 800 57922 856
rect 58090 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60590 856
rect 60758 800 60866 856
rect 61034 800 61050 856
rect 61218 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61786 856
rect 61954 800 62062 856
rect 62230 800 62246 856
rect 62414 800 62522 856
rect 62690 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63258 856
rect 63426 800 63442 856
rect 63610 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64914 856
rect 65082 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65650 856
rect 65818 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67582 856
rect 67750 800 67766 856
rect 67934 800 68042 856
rect 68210 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69238 856
rect 69406 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70250 856
rect 70418 800 70434 856
rect 70602 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71170 856
rect 71338 800 71446 856
rect 71614 800 71630 856
rect 71798 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72366 856
rect 72534 800 72642 856
rect 72810 800 72826 856
rect 72994 800 73102 856
rect 73270 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74298 856
rect 74466 800 74574 856
rect 74742 800 74758 856
rect 74926 800 75034 856
rect 75202 800 75218 856
rect 75386 800 75494 856
rect 75662 800 75770 856
rect 75938 800 75954 856
rect 76122 800 76230 856
rect 76398 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76966 856
rect 77134 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77702 856
rect 77870 800 77886 856
rect 78054 800 78162 856
rect 78330 800 78346 856
rect 78514 800 78622 856
rect 78790 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79818 856
rect 79986 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80554 856
rect 80722 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81750 856
rect 81918 800 82026 856
rect 82194 800 82210 856
rect 82378 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83406 856
rect 83574 800 83682 856
rect 83850 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84418 856
rect 84586 800 84602 856
rect 84770 800 84878 856
rect 85046 800 85154 856
rect 85322 800 85338 856
rect 85506 800 85614 856
rect 85782 800 85798 856
rect 85966 800 86074 856
rect 86242 800 86350 856
rect 86518 800 86534 856
rect 86702 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87270 856
rect 87438 800 87546 856
rect 87714 800 87730 856
rect 87898 800 88006 856
rect 88174 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89202 856
rect 89370 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89938 856
rect 90106 800 90122 856
rect 90290 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91134 856
rect 91302 800 91410 856
rect 91578 800 91594 856
rect 91762 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92606 856
rect 92774 800 92790 856
rect 92958 800 93066 856
rect 93234 800 93250 856
rect 93418 800 93526 856
rect 93694 800 93802 856
rect 93970 800 93986 856
rect 94154 800 94262 856
rect 94430 800 94446 856
rect 94614 800 94722 856
rect 94890 800 94998 856
rect 95166 800 95182 856
rect 95350 800 95458 856
rect 95626 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96654 856
rect 96822 800 96930 856
rect 97098 800 97114 856
rect 97282 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97850 856
rect 98018 800 98126 856
rect 98294 800 98310 856
rect 98478 800 98586 856
rect 98754 800 98862 856
rect 99030 800 99046 856
rect 99214 800 99322 856
rect 99490 800 99506 856
rect 99674 800 99782 856
rect 99950 800 100058 856
rect 100226 800 100242 856
rect 100410 800 100518 856
rect 100686 800 100702 856
rect 100870 800 100978 856
rect 101146 800 101254 856
rect 101422 800 101438 856
rect 101606 800 101714 856
rect 101882 800 101990 856
rect 102158 800 102174 856
rect 102342 800 102450 856
rect 102618 800 102634 856
rect 102802 800 102910 856
rect 103078 800 103186 856
rect 103354 800 103370 856
rect 103538 800 103646 856
rect 103814 800 103830 856
rect 103998 800 104106 856
rect 104274 800 104382 856
rect 104550 800 104566 856
rect 104734 800 104842 856
rect 105010 800 105026 856
rect 105194 800 105302 856
rect 105470 800 105578 856
rect 105746 800 105762 856
rect 105930 800 106038 856
rect 106206 800 106314 856
rect 106482 800 106498 856
rect 106666 800 106774 856
rect 106942 800 106958 856
rect 107126 800 107234 856
rect 107402 800 107510 856
rect 107678 800 107694 856
rect 107862 800 107970 856
rect 108138 800 108154 856
rect 108322 800 108430 856
rect 108598 800 108706 856
rect 108874 800 108890 856
rect 109058 800 109166 856
rect 109334 800 109442 856
rect 109610 800 109626 856
rect 109794 800 109902 856
rect 110070 800 110086 856
rect 110254 800 110362 856
rect 110530 800 110638 856
rect 110806 800 110822 856
rect 110990 800 111098 856
rect 111266 800 111282 856
rect 111450 800 111558 856
rect 111726 800 111834 856
rect 112002 800 112018 856
rect 112186 800 112294 856
rect 112462 800 112478 856
rect 112646 800 112754 856
rect 112922 800 113030 856
rect 113198 800 113214 856
rect 113382 800 113490 856
rect 113658 800 113766 856
rect 113934 800 113950 856
rect 114118 800 114226 856
rect 114394 800 114410 856
rect 114578 800 114686 856
rect 114854 800 114962 856
rect 115130 800 115146 856
rect 115314 800 115422 856
rect 115590 800 115606 856
rect 115774 800 115882 856
rect 116050 800 116158 856
rect 116326 800 116342 856
rect 116510 800 116618 856
rect 116786 800 116894 856
rect 117062 800 117078 856
rect 117246 800 117354 856
rect 117522 800 117538 856
rect 117706 800 117814 856
rect 117982 800 118090 856
rect 118258 800 118274 856
rect 118442 800 118478 856
<< metal3 >>
rect 0 113296 800 113416
rect 119200 113296 120000 113416
rect 0 99968 800 100088
rect 119200 99968 120000 100088
rect 0 86640 800 86760
rect 119200 86640 120000 86760
rect 0 73312 800 73432
rect 119200 73312 120000 73432
rect 0 59984 800 60104
rect 119200 59984 120000 60104
rect 0 46656 800 46776
rect 119200 46656 120000 46776
rect 0 33328 800 33448
rect 119200 33328 120000 33448
rect 0 20000 800 20120
rect 119200 20000 120000 20120
rect 0 6672 800 6792
rect 119200 6672 120000 6792
<< obsm3 >>
rect 105 113496 119200 117537
rect 880 113216 119120 113496
rect 105 100168 119200 113216
rect 880 99888 119120 100168
rect 105 86840 119200 99888
rect 880 86560 119120 86840
rect 105 73512 119200 86560
rect 880 73232 119120 73512
rect 105 60184 119200 73232
rect 880 59904 119120 60184
rect 105 46856 119200 59904
rect 880 46576 119120 46856
rect 105 33528 119200 46576
rect 880 33248 119120 33528
rect 105 20200 119200 33248
rect 880 19920 119120 20200
rect 105 6872 119200 19920
rect 880 6592 119120 6872
rect 105 1395 119200 6592
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 12203 2483 12269 3637
<< labels >>
rlabel metal2 s 115386 119200 115442 120000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 118606 0 118662 800 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 116398 119200 116454 120000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 119200 86640 120000 86760 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 118790 0 118846 800 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 0 46656 800 46776 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 119200 99968 120000 100088 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 119200 113296 120000 113416 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 117410 119200 117466 120000 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 119066 0 119122 800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 118146 0 118202 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 118422 119200 118478 120000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 119342 0 119398 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 73312 800 73432 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 119526 0 119582 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 86640 800 86760 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 119802 0 119858 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 99968 800 100088 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 119434 119200 119490 120000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 113296 800 113416 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 6672 800 6792 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal2 s 118330 0 118386 800 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 119200 33328 120000 33448 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 119200 46656 120000 46776 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 0 20000 800 20120 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 119200 59984 120000 60104 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal3 s 119200 73312 120000 73432 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 0 33328 800 33448 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 478 119200 534 120000 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 30654 119200 30710 120000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 33690 119200 33746 120000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 36726 119200 36782 120000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 39762 119200 39818 120000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 42798 119200 42854 120000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 45834 119200 45890 120000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 48778 119200 48834 120000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 51814 119200 51870 120000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 54850 119200 54906 120000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 57886 119200 57942 120000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 3422 119200 3478 120000 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 60922 119200 60978 120000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 63958 119200 64014 120000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 66994 119200 67050 120000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 70030 119200 70086 120000 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 72974 119200 73030 120000 6 io_in[24]
port 46 nsew signal input
rlabel metal2 s 76010 119200 76066 120000 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 79046 119200 79102 120000 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 82082 119200 82138 120000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 85118 119200 85174 120000 6 io_in[28]
port 50 nsew signal input
rlabel metal2 s 88154 119200 88210 120000 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 6458 119200 6514 120000 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 91190 119200 91246 120000 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 94226 119200 94282 120000 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 97170 119200 97226 120000 6 io_in[32]
port 55 nsew signal input
rlabel metal2 s 100206 119200 100262 120000 6 io_in[33]
port 56 nsew signal input
rlabel metal2 s 103242 119200 103298 120000 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 106278 119200 106334 120000 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 109314 119200 109370 120000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 9494 119200 9550 120000 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 12530 119200 12586 120000 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 15566 119200 15622 120000 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 18602 119200 18658 120000 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 21638 119200 21694 120000 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 24582 119200 24638 120000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 27618 119200 27674 120000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 31666 119200 31722 120000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 34702 119200 34758 120000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 37738 119200 37794 120000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 40774 119200 40830 120000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 43810 119200 43866 120000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 46846 119200 46902 120000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 49790 119200 49846 120000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 55862 119200 55918 120000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 58898 119200 58954 120000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 4434 119200 4490 120000 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 61934 119200 61990 120000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 64970 119200 65026 120000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 68006 119200 68062 120000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 71042 119200 71098 120000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal2 s 73986 119200 74042 120000 6 io_oeb[24]
port 84 nsew signal output
rlabel metal2 s 77022 119200 77078 120000 6 io_oeb[25]
port 85 nsew signal output
rlabel metal2 s 80058 119200 80114 120000 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 83094 119200 83150 120000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 86130 119200 86186 120000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 7470 119200 7526 120000 6 io_oeb[2]
port 90 nsew signal output
rlabel metal2 s 92202 119200 92258 120000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 95238 119200 95294 120000 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 98182 119200 98238 120000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal2 s 101218 119200 101274 120000 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 104254 119200 104310 120000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 107290 119200 107346 120000 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 110326 119200 110382 120000 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 113362 119200 113418 120000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 10506 119200 10562 120000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 13542 119200 13598 120000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 16578 119200 16634 120000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 19614 119200 19670 120000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 22650 119200 22706 120000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 25594 119200 25650 120000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 28630 119200 28686 120000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 2410 119200 2466 120000 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 32678 119200 32734 120000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 35714 119200 35770 120000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 38750 119200 38806 120000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 41786 119200 41842 120000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 44822 119200 44878 120000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 47858 119200 47914 120000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 50802 119200 50858 120000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 53838 119200 53894 120000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 56874 119200 56930 120000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 59910 119200 59966 120000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 5446 119200 5502 120000 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 62946 119200 63002 120000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 65982 119200 66038 120000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 69018 119200 69074 120000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 72054 119200 72110 120000 6 io_out[23]
port 121 nsew signal output
rlabel metal2 s 74998 119200 75054 120000 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 78034 119200 78090 120000 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 81070 119200 81126 120000 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 84106 119200 84162 120000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 87142 119200 87198 120000 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 90178 119200 90234 120000 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 8482 119200 8538 120000 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 93214 119200 93270 120000 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 io_out[31]
port 130 nsew signal output
rlabel metal2 s 99194 119200 99250 120000 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 102230 119200 102286 120000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 105266 119200 105322 120000 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 108302 119200 108358 120000 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 111338 119200 111394 120000 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 114374 119200 114430 120000 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 11518 119200 11574 120000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 14554 119200 14610 120000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 17590 119200 17646 120000 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 20626 119200 20682 120000 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 23662 119200 23718 120000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 26606 119200 26662 120000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 29642 119200 29698 120000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 user_irq[0]
port 528 nsew signal output
rlabel metal3 s 119200 6672 120000 6792 6 user_irq[1]
port 529 nsew signal output
rlabel metal3 s 119200 20000 120000 20120 6 user_irq[2]
port 530 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 531 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 531 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 531 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 531 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 532 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 532 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 532 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 532 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_ack_o
port 535 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[0]
port 601 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[10]
port 602 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[11]
port 603 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[12]
port 604 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[13]
port 605 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[14]
port 606 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[15]
port 607 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[16]
port 608 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[17]
port 609 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[18]
port 610 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[19]
port 611 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[1]
port 612 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[20]
port 613 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[21]
port 614 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[22]
port 615 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[23]
port 616 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[24]
port 617 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[25]
port 618 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[26]
port 619 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[27]
port 620 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[28]
port 621 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[29]
port 622 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[2]
port 623 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[30]
port 624 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_o[31]
port 625 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[3]
port 626 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[4]
port 627 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[5]
port 628 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[6]
port 629 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[7]
port 630 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[8]
port 631 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[9]
port 632 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4224116
string GDS_FILE /home/ren/Projects/caravel_tutorial/caravel_example/openlane/NNgen/runs/NNgen/results/finishing/basic.magic.gds
string GDS_START 173926
<< end >>

